module mspi_top
