module mspi_top
i
